module sine_lut #(
	 parameter OUTPUT_WIDTH = 12,          // 输出值位宽
	 parameter ROM_ADDR_WIDTH = 8
)(
    input wire [ROM_ADDR_WIDTH-1:0] addr,       // 8位地址
    output reg signed [OUTPUT_WIDTH-1:0] data       // 12位正弦数据
);

    always @(*) begin
        case(addr)
				 8'd0  : data = 12'sd0;
				 8'd1  : data = 12'sd50;
				 8'd2  : data = 12'sd100;
				 8'd3  : data = 12'sd151;
				 8'd4  : data = 12'sd201;
				 8'd5  : data = 12'sd251;
				 8'd6  : data = 12'sd300;
				 8'd7  : data = 12'sd350;
				 8'd8  : data = 12'sd399;
				 8'd9  : data = 12'sd449;
				 8'd10 : data = 12'sd497;
				 8'd11 : data = 12'sd546;
				 8'd12 : data = 12'sd594;
				 8'd13 : data = 12'sd642;
				 8'd14 : data = 12'sd690;
				 8'd15 : data = 12'sd737;
				 8'd16 : data = 12'sd783;
				 8'd17 : data = 12'sd830;
				 8'd18 : data = 12'sd875;
				 8'd19 : data = 12'sd920;
				 8'd20 : data = 12'sd965;
				 8'd21 : data = 12'sd1009;
				 8'd22 : data = 12'sd1052;
				 8'd23 : data = 12'sd1095;
				 8'd24 : data = 12'sd1137;
				 8'd25 : data = 12'sd1179;
				 8'd26 : data = 12'sd1219;
				 8'd27 : data = 12'sd1259;
				 8'd28 : data = 12'sd1299;
				 8'd29 : data = 12'sd1337;
				 8'd30 : data = 12'sd1375;
				 8'd31 : data = 12'sd1411;
				 8'd32 : data = 12'sd1447;
				 8'd33 : data = 12'sd1483;
				 8'd34 : data = 12'sd1517;
				 8'd35 : data = 12'sd1550;
				 8'd36 : data = 12'sd1582;
				 8'd37 : data = 12'sd1614;
				 8'd38 : data = 12'sd1644;
				 8'd39 : data = 12'sd1674;
				 8'd40 : data = 12'sd1702;
				 8'd41 : data = 12'sd1729;
				 8'd42 : data = 12'sd1756;
				 8'd43 : data = 12'sd1781;
				 8'd44 : data = 12'sd1805;
				 8'd45 : data = 12'sd1828;
				 8'd46 : data = 12'sd1850;
				 8'd47 : data = 12'sd1871;
				 8'd48 : data = 12'sd1891;
				 8'd49 : data = 12'sd1910;
				 8'd50 : data = 12'sd1927;
				 8'd51 : data = 12'sd1944;
				 8'd52 : data = 12'sd1959;
				 8'd53 : data = 12'sd1973;
				 8'd54 : data = 12'sd1986;
				 8'd55 : data = 12'sd1997;
				 8'd56 : data = 12'sd2008;
				 8'd57 : data = 12'sd2017;
				 8'd58 : data = 12'sd2025;
				 8'd59 : data = 12'sd2032;
				 8'd60 : data = 12'sd2037;
				 8'd61 : data = 12'sd2041;
				 8'd62 : data = 12'sd2045;
				 8'd63 : data = 12'sd2046;
				 8'd64 : data = 12'sd2047;
				 8'd65 : data = 12'sd2046;
				 8'd66 : data = 12'sd2045;
				 8'd67 : data = 12'sd2041;
				 8'd68 : data = 12'sd2037;
				 8'd69 : data = 12'sd2032;
				 8'd70 : data = 12'sd2025;
				 8'd71 : data = 12'sd2017;
				 8'd72 : data = 12'sd2008;
				 8'd73 : data = 12'sd1997;
				 8'd74 : data = 12'sd1986;
				 8'd75 : data = 12'sd1973;
				 8'd76 : data = 12'sd1959;
				 8'd77 : data = 12'sd1944;
				 8'd78 : data = 12'sd1927;
				 8'd79 : data = 12'sd1910;
				 8'd80 : data = 12'sd1891;
				 8'd81 : data = 12'sd1871;
				 8'd82 : data = 12'sd1850;
				 8'd83 : data = 12'sd1828;
				 8'd84 : data = 12'sd1805;
				 8'd85 : data = 12'sd1781;
				 8'd86 : data = 12'sd1756;
				 8'd87 : data = 12'sd1729;
				 8'd88 : data = 12'sd1702;
				 8'd89 : data = 12'sd1674;
				 8'd90 : data = 12'sd1644;
				 8'd91 : data = 12'sd1614;
				 8'd92 : data = 12'sd1582;
				 8'd93 : data = 12'sd1550;
				 8'd94 : data = 12'sd1517;
				 8'd95 : data = 12'sd1483;
				 8'd96 : data = 12'sd1447;
				 8'd97 : data = 12'sd1411;
				 8'd98 : data = 12'sd1375;
				 8'd99 : data = 12'sd1337;
				 8'd100: data = 12'sd1299;
				 8'd101: data = 12'sd1259;
				 8'd102: data = 12'sd1219;
				 8'd103: data = 12'sd1179;
				 8'd104: data = 12'sd1137;
				 8'd105: data = 12'sd1095;
				 8'd106: data = 12'sd1052;
				 8'd107: data = 12'sd1009;
				 8'd108: data = 12'sd965;
				 8'd109: data = 12'sd920;
				 8'd110: data = 12'sd875;
				 8'd111: data = 12'sd830;
				 8'd112: data = 12'sd783;
				 8'd113: data = 12'sd737;
				 8'd114: data = 12'sd690;
				 8'd115: data = 12'sd642;
				 8'd116: data = 12'sd594;
				 8'd117: data = 12'sd546;
				 8'd118: data = 12'sd497;
				 8'd119: data = 12'sd449;
				 8'd120: data = 12'sd399;
				 8'd121: data = 12'sd350;
				 8'd122: data = 12'sd300;
				 8'd123: data = 12'sd251;
				 8'd124: data = 12'sd201;
				 8'd125: data = 12'sd151;
				 8'd126: data = 12'sd100;
				 8'd127: data = 12'sd50;
				 8'd128: data = 12'sd0;
				 8'd129: data = -12'sd50;
				 8'd130: data = -12'sd100;
				 8'd131: data = -12'sd151;
				 8'd132: data = -12'sd201;
				 8'd133: data = -12'sd251;
				 8'd134: data = -12'sd300;
				 8'd135: data = -12'sd350;
				 8'd136: data = -12'sd399;
				 8'd137: data = -12'sd449;
				 8'd138: data = -12'sd497;
				 8'd139: data = -12'sd546;
				 8'd140: data = -12'sd594;
				 8'd141: data = -12'sd642;
				 8'd142: data = -12'sd690;
				 8'd143: data = -12'sd737;
				 8'd144: data = -12'sd783;
				 8'd145: data = -12'sd830;
				 8'd146: data = -12'sd875;
				 8'd147: data = -12'sd920;
				 8'd148: data = -12'sd965;
				 8'd149: data = -12'sd1009;
				 8'd150: data = -12'sd1052;
				 8'd151: data = -12'sd1095;
				 8'd152: data = -12'sd1137;
				 8'd153: data = -12'sd1179;
				 8'd154: data = -12'sd1219;
				 8'd155: data = -12'sd1259;
				 8'd156: data = -12'sd1299;
				 8'd157: data = -12'sd1337;
				 8'd158: data = -12'sd1375;
				 8'd159: data = -12'sd1411;
				 8'd160: data = -12'sd1447;
				 8'd161: data = -12'sd1483;
				 8'd162: data = -12'sd1517;
				 8'd163: data = -12'sd1550;
				 8'd164: data = -12'sd1582;
				 8'd165: data = -12'sd1614;
				 8'd166: data = -12'sd1644;
				 8'd167: data = -12'sd1674;
				 8'd168: data = -12'sd1702;
				 8'd169: data = -12'sd1729;
				 8'd170: data = -12'sd1756;
				 8'd171: data = -12'sd1781;
				 8'd172: data = -12'sd1805;
				 8'd173: data = -12'sd1828;
				 8'd174: data = -12'sd1850;
				 8'd175: data = -12'sd1871;
				 8'd176: data = -12'sd1891;
				 8'd177: data = -12'sd1910;
				 8'd178: data = -12'sd1927;
				 8'd179: data = -12'sd1944;
				 8'd180: data = -12'sd1959;
				 8'd181: data = -12'sd1973;
				 8'd182: data = -12'sd1986;
				 8'd183: data = -12'sd1997;
				 8'd184: data = -12'sd2008;
				 8'd185: data = -12'sd2017;
				 8'd186: data = -12'sd2025;
				 8'd187: data = -12'sd2032;
				 8'd188: data = -12'sd2037;
				 8'd189: data = -12'sd2041;
				 8'd190: data = -12'sd2045;
				 8'd191: data = -12'sd2046;
				 8'd192: data = -12'sd2047;
				 8'd193: data = -12'sd2046;
				 8'd194: data = -12'sd2045;
				 8'd195: data = -12'sd2041;
				 8'd196: data = -12'sd2037;
				 8'd197: data = -12'sd2032;
				 8'd198: data = -12'sd2025;
				 8'd199: data = -12'sd2017;
				 8'd200: data = -12'sd2008;
				 8'd201: data = -12'sd1997;
				 8'd202: data = -12'sd1986;
				 8'd203: data = -12'sd1973;
				 8'd204: data = -12'sd1959;
				 8'd205: data = -12'sd1944;
				 8'd206: data = -12'sd1927;
				 8'd207: data = -12'sd1910;
				 8'd208: data = -12'sd1891;
				 8'd209: data = -12'sd1871;
				 8'd210: data = -12'sd1850;
				 8'd211: data = -12'sd1828;
				 8'd212: data = -12'sd1805;
				 8'd213: data = -12'sd1781;
				 8'd214: data = -12'sd1756;
				 8'd215: data = -12'sd1729;
				 8'd216: data = -12'sd1702;
				 8'd217: data = -12'sd1674;
				 8'd218: data = -12'sd1644;
				 8'd219: data = -12'sd1614;
				 8'd220: data = -12'sd1582;
				 8'd221: data = -12'sd1550;
				 8'd222: data = -12'sd1517;
				 8'd223: data = -12'sd1483;
				 8'd224: data = -12'sd1447;
				 8'd225: data = -12'sd1411;
				 8'd226: data = -12'sd1375;
				 8'd227: data = -12'sd1337;
				 8'd228: data = -12'sd1299;
				 8'd229: data = -12'sd1259;
				 8'd230: data = -12'sd1219;
				 8'd231: data = -12'sd1179;
				 8'd232: data = -12'sd1137;
				 8'd233: data = -12'sd1095;
				 8'd234: data = -12'sd1052;
				 8'd235: data = -12'sd1009;
				 8'd236: data = -12'sd965;
				 8'd237: data = -12'sd920;
				 8'd238: data = -12'sd875;
				 8'd239: data = -12'sd830;
				 8'd240: data = -12'sd783;
				 8'd241: data = -12'sd737;
				 8'd242: data = -12'sd690;
				 8'd243: data = -12'sd642;
				 8'd244: data = -12'sd594;
				 8'd245: data = -12'sd546;
				 8'd246: data = -12'sd497;
				 8'd247: data = -12'sd449;
				 8'd248: data = -12'sd399;
				 8'd249: data = -12'sd350;
				 8'd250: data = -12'sd300;
				 8'd251: data = -12'sd251;
				 8'd252: data = -12'sd201;
				 8'd253: data = -12'sd151;
				 8'd254: data = -12'sd100;
				 8'd255: data = -12'sd50;
			endcase
    end

endmodule