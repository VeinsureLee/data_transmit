module sine_lut #(
	 parameter OUTPUT_WIDTH = 12,          // 输出值位宽
	 parameter ROM_ADDR_WIDTH = 8
)(
    input wire [ROM_ADDR_WIDTH-1:0] addr,       // 8位地址
    output reg [OUTPUT_WIDTH-1:0] data       // 12位正弦数据
);

    always @(*) begin
        case(addr)
            8'd0:   data = 12'd2048;
            8'd1:   data = 12'd2073;
            8'd2:   data = 12'd2097;
            8'd3:   data = 12'd2122;
            8'd4:   data = 12'd2146;
            8'd5:   data = 12'd2170;
            8'd6:   data = 12'd2195;
            8'd7:   data = 12'd2219;
            8'd8:   data = 12'd2243;
            8'd9:   data = 12'd2267;
            8'd10:   data = 12'd2291;
            8'd11:   data = 12'd2315;
            8'd12:   data = 12'd2338;
            8'd13:   data = 12'd2362;
            8'd14:   data = 12'd2385;
            8'd15:   data = 12'd2408;
            8'd16:   data = 12'd2431;
            8'd17:   data = 12'd2453;
            8'd18:   data = 12'd2476;
            8'd19:   data = 12'd2498;
            8'd20:   data = 12'd2519;
            8'd21:   data = 12'd2541;
            8'd22:   data = 12'd2562;
            8'd23:   data = 12'd2583;
            8'd24:   data = 12'd2604;
            8'd25:   data = 12'd2624;
            8'd26:   data = 12'd2644;
            8'd27:   data = 12'd2663;
            8'd28:   data = 12'd2682;
            8'd29:   data = 12'd2701;
            8'd30:   data = 12'd2720;
            8'd31:   data = 12'd2738;
            8'd32:   data = 12'd2755;
            8'd33:   data = 12'd2772;
            8'd34:   data = 12'd2789;
            8'd35:   data = 12'd2805;
            8'd36:   data = 12'd2821;
            8'd37:   data = 12'd2836;
            8'd38:   data = 12'd2851;
            8'd39:   data = 12'd2866;
            8'd40:   data = 12'd2879;
            8'd41:   data = 12'd2893;
            8'd42:   data = 12'd2906;
            8'd43:   data = 12'd2918;
            8'd44:   data = 12'd2930;
            8'd45:   data = 12'd2941;
            8'd46:   data = 12'd2952;
            8'd47:   data = 12'd2962;
            8'd48:   data = 12'd2972;
            8'd49:   data = 12'd2981;
            8'd50:   data = 12'd2990;
            8'd51:   data = 12'd2998;
            8'd52:   data = 12'd3005;
            8'd53:   data = 12'd3012;
            8'd54:   data = 12'd3018;
            8'd55:   data = 12'd3024;
            8'd56:   data = 12'd3029;
            8'd57:   data = 12'd3033;
            8'd58:   data = 12'd3037;
            8'd59:   data = 12'd3040;
            8'd60:   data = 12'd3043;
            8'd61:   data = 12'd3045;
            8'd62:   data = 12'd3047;
            8'd63:   data = 12'd3048;
            8'd64:   data = 12'd3048;
            8'd65:   data = 12'd3048;
            8'd66:   data = 12'd3047;
            8'd67:   data = 12'd3045;
            8'd68:   data = 12'd3043;
            8'd69:   data = 12'd3040;
            8'd70:   data = 12'd3037;
            8'd71:   data = 12'd3033;
            8'd72:   data = 12'd3029;
            8'd73:   data = 12'd3024;
            8'd74:   data = 12'd3018;
            8'd75:   data = 12'd3012;
            8'd76:   data = 12'd3005;
            8'd77:   data = 12'd2998;
            8'd78:   data = 12'd2990;
            8'd79:   data = 12'd2981;
            8'd80:   data = 12'd2972;
            8'd81:   data = 12'd2962;
            8'd82:   data = 12'd2952;
            8'd83:   data = 12'd2941;
            8'd84:   data = 12'd2930;
            8'd85:   data = 12'd2918;
            8'd86:   data = 12'd2906;
            8'd87:   data = 12'd2893;
            8'd88:   data = 12'd2879;
            8'd89:   data = 12'd2866;
            8'd90:   data = 12'd2851;
            8'd91:   data = 12'd2836;
            8'd92:   data = 12'd2821;
            8'd93:   data = 12'd2805;
            8'd94:   data = 12'd2789;
            8'd95:   data = 12'd2772;
            8'd96:   data = 12'd2755;
            8'd97:   data = 12'd2738;
            8'd98:   data = 12'd2720;
            8'd99:   data = 12'd2701;
            8'd100:   data = 12'd2682;
            8'd101:   data = 12'd2663;
            8'd102:   data = 12'd2644;
            8'd103:   data = 12'd2624;
            8'd104:   data = 12'd2604;
            8'd105:   data = 12'd2583;
            8'd106:   data = 12'd2562;
            8'd107:   data = 12'd2541;
            8'd108:   data = 12'd2519;
            8'd109:   data = 12'd2498;
            8'd110:   data = 12'd2476;
            8'd111:   data = 12'd2453;
            8'd112:   data = 12'd2431;
            8'd113:   data = 12'd2408;
            8'd114:   data = 12'd2385;
            8'd115:   data = 12'd2362;
            8'd116:   data = 12'd2338;
            8'd117:   data = 12'd2315;
            8'd118:   data = 12'd2291;
            8'd119:   data = 12'd2267;
            8'd120:   data = 12'd2243;
            8'd121:   data = 12'd2219;
            8'd122:   data = 12'd2195;
            8'd123:   data = 12'd2170;
            8'd124:   data = 12'd2146;
            8'd125:   data = 12'd2122;
            8'd126:   data = 12'd2097;
            8'd127:   data = 12'd2073;
            8'd128:   data = 12'd2048;
            8'd129:   data = 12'd2023;
            8'd130:   data = 12'd1999;
            8'd131:   data = 12'd1974;
            8'd132:   data = 12'd1950;
            8'd133:   data = 12'd1926;
            8'd134:   data = 12'd1901;
            8'd135:   data = 12'd1877;
            8'd136:   data = 12'd1853;
            8'd137:   data = 12'd1829;
            8'd138:   data = 12'd1805;
            8'd139:   data = 12'd1781;
            8'd140:   data = 12'd1758;
            8'd141:   data = 12'd1734;
            8'd142:   data = 12'd1711;
            8'd143:   data = 12'd1688;
            8'd144:   data = 12'd1665;
            8'd145:   data = 12'd1643;
            8'd146:   data = 12'd1620;
            8'd147:   data = 12'd1598;
            8'd148:   data = 12'd1577;
            8'd149:   data = 12'd1555;
            8'd150:   data = 12'd1534;
            8'd151:   data = 12'd1513;
            8'd152:   data = 12'd1492;
            8'd153:   data = 12'd1472;
            8'd154:   data = 12'd1452;
            8'd155:   data = 12'd1433;
            8'd156:   data = 12'd1414;
            8'd157:   data = 12'd1395;
            8'd158:   data = 12'd1376;
            8'd159:   data = 12'd1358;
            8'd160:   data = 12'd1341;
            8'd161:   data = 12'd1324;
            8'd162:   data = 12'd1307;
            8'd163:   data = 12'd1291;
            8'd164:   data = 12'd1275;
            8'd165:   data = 12'd1260;
            8'd166:   data = 12'd1245;
            8'd167:   data = 12'd1230;
            8'd168:   data = 12'd1217;
            8'd169:   data = 12'd1203;
            8'd170:   data = 12'd1190;
            8'd171:   data = 12'd1178;
            8'd172:   data = 12'd1166;
            8'd173:   data = 12'd1155;
            8'd174:   data = 12'd1144;
            8'd175:   data = 12'd1134;
            8'd176:   data = 12'd1124;
            8'd177:   data = 12'd1115;
            8'd178:   data = 12'd1106;
            8'd179:   data = 12'd1098;
            8'd180:   data = 12'd1091;
            8'd181:   data = 12'd1084;
            8'd182:   data = 12'd1078;
            8'd183:   data = 12'd1072;
            8'd184:   data = 12'd1067;
            8'd185:   data = 12'd1063;
            8'd186:   data = 12'd1059;
            8'd187:   data = 12'd1056;
            8'd188:   data = 12'd1053;
            8'd189:   data = 12'd1051;
            8'd190:   data = 12'd1049;
            8'd191:   data = 12'd1048;
            8'd192:   data = 12'd1048;
            8'd193:   data = 12'd1048;
            8'd194:   data = 12'd1049;
            8'd195:   data = 12'd1051;
            8'd196:   data = 12'd1053;
            8'd197:   data = 12'd1056;
            8'd198:   data = 12'd1059;
            8'd199:   data = 12'd1063;
            8'd200:   data = 12'd1067;
            8'd201:   data = 12'd1072;
            8'd202:   data = 12'd1078;
            8'd203:   data = 12'd1084;
            8'd204:   data = 12'd1091;
            8'd205:   data = 12'd1098;
            8'd206:   data = 12'd1106;
            8'd207:   data = 12'd1115;
            8'd208:   data = 12'd1124;
            8'd209:   data = 12'd1134;
            8'd210:   data = 12'd1144;
            8'd211:   data = 12'd1155;
            8'd212:   data = 12'd1166;
            8'd213:   data = 12'd1178;
            8'd214:   data = 12'd1190;
            8'd215:   data = 12'd1203;
            8'd216:   data = 12'd1217;
            8'd217:   data = 12'd1230;
            8'd218:   data = 12'd1245;
            8'd219:   data = 12'd1260;
            8'd220:   data = 12'd1275;
            8'd221:   data = 12'd1291;
            8'd222:   data = 12'd1307;
            8'd223:   data = 12'd1324;
            8'd224:   data = 12'd1341;
            8'd225:   data = 12'd1358;
            8'd226:   data = 12'd1376;
            8'd227:   data = 12'd1395;
            8'd228:   data = 12'd1414;
            8'd229:   data = 12'd1433;
            8'd230:   data = 12'd1452;
            8'd231:   data = 12'd1472;
            8'd232:   data = 12'd1492;
            8'd233:   data = 12'd1513;
            8'd234:   data = 12'd1534;
            8'd235:   data = 12'd1555;
            8'd236:   data = 12'd1577;
            8'd237:   data = 12'd1598;
            8'd238:   data = 12'd1620;
            8'd239:   data = 12'd1643;
            8'd240:   data = 12'd1665;
            8'd241:   data = 12'd1688;
            8'd242:   data = 12'd1711;
            8'd243:   data = 12'd1734;
            8'd244:   data = 12'd1758;
            8'd245:   data = 12'd1781;
            8'd246:   data = 12'd1805;
            8'd247:   data = 12'd1829;
            8'd248:   data = 12'd1853;
            8'd249:   data = 12'd1877;
            8'd250:   data = 12'd1901;
            8'd251:   data = 12'd1926;
            8'd252:   data = 12'd1950;
            8'd253:   data = 12'd1974;
            8'd254:   data = 12'd1999;
            8'd255:   data = 12'd2023;
            default: data = 12'd2048;
        endcase
    end

endmodule
